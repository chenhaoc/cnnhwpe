`define D_Kernel_size 11
`define D_Data_type 3
`define D_Layer_type 1
`define D_Kernel_333 0
`define D_H 25
`define D_W 25
`define D_C 3
`define D_K 32
`define D_STRIDE 2
`define D_fmap_file_path ".\\case_gen_txt\\conv_input_11str2\\inputimage_11.bin"
`define D_kernel_file_path ".\\case_gen_txt\\conv_input_11str2\\inputfilter_11.bin"
`define D_conv_file_path ".\\case_gen_txt\\conv_input_11str2\\conv_11.bin"
