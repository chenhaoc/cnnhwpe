`define D_Kernel_size 3
`define D_Data_type 2
`define D_Layer_type 0
`define D_Kernel_333 0
`define D_H 17
`define D_W 17
`define D_C 32
`define D_K 32
`define D_STRIDE 2
`define D_fmap_file_path ".\\case_gen_txt\\conv_input_4bstr2\\featuremap_4b.bin"
`define D_kernel_file_path ".\\case_gen_txt\\conv_input_4bstr2\\fmapfilter_4b.bin"
`define D_conv_file_path ".\\case_gen_txt\\conv_input_4bstr2\\conv_4b.bin"
