`define D_Kernel_size 3
`define D_Data_type 3
`define D_Layer_type 0
`define D_Kernel_333 0
`define D_H 10
`define D_W 10
`define D_C 32
`define D_K 32
`define D_STRIDE 1
`define D_fmap_file_path ".\\case_gen_txt\\conv_input_3str1\\featuremap_8b.bin"
`define D_kernel_file_path ".\\case_gen_txt\\conv_input_3str1\\fmapfilter_8b.bin"
`define D_conv_file_path ".\\case_gen_txt\\conv_input_3str1\\conv_8b.bin"
