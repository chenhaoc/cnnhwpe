`define D_Kernel_size 3
`define D_Data_type 3
`define D_Layer_type 1
`define D_Kernel_333 1
`define D_H 10
`define D_W 10
`define D_C 3
`define D_K 32
`define D_STRIDE 1
`define D_fmap_file_path ".\\case_gen_txt\\conv_input_3str1\\inputimage_3.bin"
`define D_kernel_file_path ".\\case_gen_txt\\conv_input_3str1\\inputfilter_3.bin"
`define D_conv_file_path ".\\case_gen_txt\\conv_input_3str1\\conv_3.bin"
